../08_dev_loader/dev_io_switch.sv