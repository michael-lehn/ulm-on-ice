../10_io_interface/uart_tx.sv