../11_ram/dev_ram.sv