../13_ram32/if_ram.sv