../13_ram32/dev_ram.sv