../08_dev_loader/dev_ram.sv