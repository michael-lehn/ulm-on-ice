../13_ram32/long_we_mask.sv