../07_io_interface/fifo.sv