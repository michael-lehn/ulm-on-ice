../07_io_interface/pkg_ram.sv