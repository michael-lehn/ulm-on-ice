../11_ram/SB_SPRAM256KA.sv