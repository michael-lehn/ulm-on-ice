../06_io_mirror/baud_tick_gen.sv