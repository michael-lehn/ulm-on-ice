interface if_iobuf;
    logic empty;
    logic [7:0] data_out;
    logic pop_front;
    logic full;
    logic push_back;
    logic [7:0] data_in;
endinterface

