../08_dev_loader/SB_SPRAM256KA.sv