../08_dev_loader/dev_loader.sv