../13_ram32/long_ext_high.sv