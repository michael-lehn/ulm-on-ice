../10_io_interface/fifo.sv