../13_ram32/long_rshift.sv