../11_ram/pkg_ram.sv