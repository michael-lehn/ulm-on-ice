../11_ram/quad_rshift.sv