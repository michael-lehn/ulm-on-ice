../07_io_interface/dev_hex.sv