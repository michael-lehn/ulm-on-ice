../08_dev_loader/if_ram.sv