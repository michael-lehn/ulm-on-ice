../13_ram32/spram.sv