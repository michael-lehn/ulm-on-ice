../08_dev_loader/quad_lshift.sv