../11_ram/quad_ext_low.sv