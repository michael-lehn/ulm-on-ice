../07_io_interface/dp_bram4096.sv