../11_ram/if_ram.sv