../03_hexdisplay/dev_hex.sv