../08_dev_loader/quad_we_mask.sv