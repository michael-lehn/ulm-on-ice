../11_ram/quad_ext_high.sv