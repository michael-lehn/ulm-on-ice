../04_dip_switch/dev_hex.sv