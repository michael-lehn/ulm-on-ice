../07_io_interface/if_fifo.sv