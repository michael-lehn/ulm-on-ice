../11_ram/spram.sv