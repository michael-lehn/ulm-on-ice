../13_ram32/pkg_ram.sv