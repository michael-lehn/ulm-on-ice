../07_io_interface/dev_io.sv