../13_ram32/SB_SPRAM256KA.sv