../08_dev_loader/spram.sv