../11_ram/quad_we_mask.sv