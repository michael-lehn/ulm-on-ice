../07_io_interface/baud_tick_gen.sv