../08_dev_loader/quad_rshift.sv