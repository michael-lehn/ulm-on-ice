../11_ram/quad_lshift.sv