../08_dev_loader/dev_ram_switch.sv