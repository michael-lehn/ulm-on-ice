../10_io_interface/if_io.sv