../07_io_interface/uart_rx.sv