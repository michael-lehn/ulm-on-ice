../13_ram32/long_ext_low.sv