../13_ram32/long_lshift.sv