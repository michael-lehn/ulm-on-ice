../08_dev_loader/quad_ext_low.sv